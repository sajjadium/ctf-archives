`INSTR(ARITH,     7'b0110011, R, ALU)
`INSTR(ARITH_IMM, 7'b0010011, I, ALU) 
`INSTR(LUI,       7'b0110111, U, ALU)

`INSTR(BRANCH,    7'b1100011, B, BU)
`INSTR(JAL,       7'b1101111, J, BU)
`INSTR(JALR,      7'b1100111, I, BU)

`INSTR(LOAD,      7'b0000011, I, LSU)
`INSTR(STORE,     7'b0100011, S, LSU)

`INSTR(AUIPC,     7'b0010111, U, BU)
`INSTR(ECALL,     7'b1110011, I, BU)
`INSTR(ERET,      7'b1110010, J, BU)

`INSTR(SETPRIV,      7'b0110100, R, PU)

`INSTR(FLAG,      7'b1110000, U, IOU)
`INSTR(WELCOME,      7'b1110001, U, IOU)