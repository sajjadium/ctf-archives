module logick(CLK, RESET_N, BYTE, GOOD);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  input [7:0] BYTE;
  input CLK;
  output GOOD;
  input RESET_N;
  reg [26:0] state;
  assign _171_ = ~BYTE[0];
  assign _172_ = BYTE[1] | _171_;
  assign _173_ = ~BYTE[3];
  assign _174_ = ~(BYTE[2] & _173_);
  assign _175_ = _174_ | _172_;
  assign _176_ = BYTE[4] & BYTE[5];
  assign _177_ = ~BYTE[7];
  assign _178_ = _177_ & BYTE[6];
  assign _179_ = ~(_178_ & _176_);
  assign _180_ = _179_ | _175_;
  assign _181_ = ~(_180_ & RESET_N);
  assign _182_ = BYTE[2] | _173_;
  assign _183_ = _182_ | _172_;
  assign _184_ = ~((_183_ | _179_) & state[1]);
  assign _185_ = ~BYTE[5];
  assign _186_ = BYTE[4] & _185_;
  assign _187_ = ~(_186_ & _178_);
  assign _188_ = BYTE[2] & BYTE[3];
  assign _189_ = BYTE[1] & BYTE[0];
  assign _190_ = ~(_189_ & _188_);
  assign _191_ = ~((_190_ | _187_) & (state[9] | state[15]));
  assign _192_ = ~((_191_ & _184_) | _181_);
  assign _193_ = ~state[22];
  assign _194_ = ~(BYTE[1] | BYTE[0]);
  assign _195_ = ~(BYTE[2] | BYTE[3]);
  assign _196_ = _195_ & _194_;
  assign _197_ = ~(BYTE[7] | BYTE[6]);
  assign _198_ = _197_ & _176_;
  assign _199_ = _198_ & _196_;
  assign _200_ = _199_ | _193_;
  assign _201_ = ~state[5];
  assign _202_ = ~(BYTE[4] | _185_);
  assign _203_ = _202_ & _178_;
  assign _204_ = BYTE[2] & _173_;
  assign _205_ = _189_ & _204_;
  assign _206_ = _205_ & _203_;
  assign _000_ = _206_ | _201_;
  assign _001_ = ~((_000_ & _200_) | _181_);
  assign _002_ = _001_ | _192_;
  assign _003_ = ~(_202_ & _178_);
  assign _004_ = _003_ | _183_;
  assign _005_ = ~(_004_ & RESET_N);
  assign _006_ = _195_ & _189_;
  assign _007_ = _006_ & _203_;
  assign _008_ = ~(_180_ & state[21]);
  assign _009_ = _008_ | _007_;
  assign _010_ = ~(_009_ | _005_);
  assign _011_ = _194_ & _188_;
  assign _012_ = _011_ & _203_;
  assign _013_ = state[8] | state[26];
  assign _014_ = ~(_013_ | state[3]);
  assign _015_ = _014_ | _012_;
  assign _016_ = ~((_015_ | _181_) & RESET_N);
  assign _017_ = _016_ | _010_;
  assign _018_ = _017_ | _002_;
  assign _019_ = ~state[7];
  assign _020_ = ~(state[0] | state[10]);
  assign _021_ = _020_ & _019_;
  assign _022_ = ~state[13];
  assign _023_ = _006_ & _198_;
  assign _024_ = _023_ | _022_;
  assign _025_ = ~((_024_ & _021_) | _181_);
  assign _026_ = ~RESET_N;
  assign _027_ = ~(_194_ & _204_);
  assign _028_ = ~(_027_ | _179_);
  assign _029_ = _028_ | _026_;
  assign _030_ = ~((state[2] | state[4]) & _180_);
  assign _031_ = BYTE[1] & _171_;
  assign _032_ = ~(_031_ & _195_);
  assign _033_ = ~((_032_ | _179_) & state[20]);
  assign _034_ = ~((_033_ | _181_) & (_030_ | _029_));
  assign _035_ = _034_ | _025_;
  assign _036_ = ~(BYTE[4] | BYTE[5]);
  assign _037_ = ~(_036_ & _178_);
  assign _038_ = ~((_037_ | _183_) & state[19]);
  assign _039_ = ~state[12];
  assign _040_ = _007_ | _039_;
  assign _041_ = ~((_040_ & _038_) | _181_);
  assign _042_ = ~(BYTE[1] | _171_);
  assign _043_ = _195_ & _042_;
  assign _044_ = ~(_043_ & _203_);
  assign _045_ = ~(_044_ & state[25]);
  assign _046_ = _178_ & _176_;
  assign _047_ = _188_ & _042_;
  assign _048_ = ~(_047_ & _046_);
  assign _049_ = ~(_048_ & state[17]);
  assign _050_ = ~((_049_ & _045_) | _181_);
  assign _051_ = _050_ | _041_;
  assign _052_ = _051_ | _035_;
  assign _053_ = _043_ & _198_;
  assign _054_ = _053_ | _026_;
  assign _055_ = ~(_180_ & state[24]);
  assign _056_ = _004_ & RESET_N;
  assign _057_ = _180_ & state[14];
  assign _058_ = _006_ & _046_;
  assign _059_ = ~(_058_ | _026_);
  assign _060_ = _180_ & state[16];
  assign _061_ = ~((_060_ & _059_) | (_057_ & _056_));
  assign _062_ = ~((_055_ | _054_) & _061_);
  assign _063_ = _031_ & _204_;
  assign _064_ = _063_ & _203_;
  assign _065_ = _064_ | _026_;
  assign _066_ = ~(_180_ & state[18]);
  assign _067_ = ~((_187_ | _175_) & state[6]);
  assign _068_ = ~((_067_ | _181_) & (_066_ | _065_));
  assign _069_ = ~(BYTE[1] & BYTE[0]);
  assign _070_ = _069_ | _182_;
  assign _071_ = ~(_070_ | _179_);
  assign _072_ = _071_ | _026_;
  assign _073_ = ~(_180_ & state[11]);
  assign _074_ = _196_ & _046_;
  assign _075_ = _074_ | _026_;
  assign _076_ = ~(_180_ & state[23]);
  assign _077_ = ~((_076_ | _075_) & (_073_ | _072_));
  assign _078_ = _077_ | _068_;
  assign _079_ = _078_ | _062_;
  assign _080_ = _079_ | _052_;
  assign _086_ = _080_ | _018_;
  assign _081_ = ~state[21];
  assign _082_ = _180_ | _081_;
  assign _083_ = _082_ | _007_;
  assign _084_ = _180_ | _026_;
  assign _085_ = ~((_049_ & _020_) | _084_);
  assign _087_ = ~((_045_ & _040_) | _084_);
  assign _088_ = ~(_087_ | _085_);
  assign _089_ = ~((_083_ | _005_) & _088_);
  assign _090_ = ~((_015_ & _184_) | _084_);
  assign _091_ = ~((_033_ & _024_) | _084_);
  assign _092_ = _091_ | _090_;
  assign _093_ = ~((_038_ & _000_) | _084_);
  assign _094_ = ~((_200_ & _191_) | _084_);
  assign _095_ = _094_ | _093_;
  assign _096_ = _095_ | _092_;
  assign _097_ = ~state[11];
  assign _098_ = _180_ | _097_;
  assign _099_ = ~state[18];
  assign _100_ = _180_ | _099_;
  assign _101_ = ~((_100_ | _065_) & (_098_ | _072_));
  assign _102_ = ~(state[2] | state[4]);
  assign _103_ = _102_ | _180_;
  assign _104_ = ~state[14];
  assign _105_ = _180_ | _104_;
  assign _106_ = ~((_105_ | _005_) & (_103_ | _029_));
  assign _107_ = _106_ | _101_;
  assign _108_ = ~state[23];
  assign _109_ = _180_ | _108_;
  assign _110_ = ~((_109_ | _075_) & (_084_ | _067_));
  assign _111_ = _058_ | _026_;
  assign _112_ = ~state[16];
  assign _113_ = _180_ | _112_;
  assign _114_ = ~state[24];
  assign _115_ = _180_ | _114_;
  assign _116_ = ~((_115_ | _054_) & (_113_ | _111_));
  assign _117_ = _116_ | _110_;
  assign _118_ = _117_ | _107_;
  assign _119_ = _118_ | _096_;
  assign _135_ = _119_ | _089_;
  assign _120_ = _004_ | _026_;
  assign _121_ = _007_ | _081_;
  assign _142_ = ~((_121_ & _104_) | _120_);
  assign _122_ = ~(state[25] & RESET_N);
  assign _147_ = ~(_122_ | _044_);
  assign _123_ = _007_ & RESET_N;
  assign _148_ = _123_ & state[21];
  assign _124_ = state[22] & RESET_N;
  assign _149_ = _124_ & _199_;
  assign _125_ = state[23] & RESET_N;
  assign _150_ = _125_ & _074_;
  assign _126_ = ~(_183_ | _179_);
  assign _127_ = state[1] & RESET_N;
  assign _151_ = _127_ & _126_;
  assign _128_ = _012_ & RESET_N;
  assign _152_ = _128_ & state[3];
  assign _129_ = ~(_187_ | _175_);
  assign _130_ = state[6] & RESET_N;
  assign _153_ = _130_ & _129_;
  assign _154_ = _123_ & state[12];
  assign _131_ = ~(state[17] & RESET_N);
  assign _155_ = ~(_131_ | _048_);
  assign _132_ = state[24] & RESET_N;
  assign _156_ = _132_ & _053_;
  assign _133_ = state[18] & RESET_N;
  assign _157_ = _133_ & _064_;
  assign _158_ = _128_ & state[26];
  assign _134_ = _028_ & RESET_N;
  assign _159_ = _134_ & state[2];
  assign _160_ = _134_ & state[4];
  assign _136_ = state[5] & RESET_N;
  assign _161_ = _136_ & _206_;
  assign _162_ = ~(_084_ | _019_);
  assign _163_ = _128_ & state[8];
  assign _137_ = ~(_190_ | _187_);
  assign _138_ = _137_ & RESET_N;
  assign _164_ = _138_ & state[9];
  assign _139_ = state[11] & RESET_N;
  assign _165_ = _139_ & _071_;
  assign _140_ = state[13] & RESET_N;
  assign _166_ = _140_ & _023_;
  assign _167_ = _138_ & state[15];
  assign _141_ = state[16] & RESET_N;
  assign _168_ = _141_ & _058_;
  assign _143_ = ~(_037_ | _183_);
  assign _144_ = state[19] & RESET_N;
  assign _169_ = _144_ & _143_;
  assign _145_ = ~(_032_ | _179_);
  assign _146_ = state[20] & RESET_N;
  assign _170_ = _146_ & _145_;
  always @(posedge CLK)
      state[0] <= _086_;
  always @(posedge CLK)
      state[1] <= _158_;
  always @(posedge CLK)
      state[2] <= _156_;
  always @(posedge CLK)
      state[3] <= _147_;
  always @(posedge CLK)
      state[4] <= _148_;
  always @(posedge CLK)
      state[5] <= _149_;
  always @(posedge CLK)
      state[6] <= _150_;
  always @(posedge CLK)
      state[7] <= _142_;
  always @(posedge CLK)
      state[8] <= _167_;
  always @(posedge CLK)
      state[9] <= _168_;
  always @(posedge CLK)
      state[10] <= _155_;
  always @(posedge CLK)
      state[11] <= _157_;
  always @(posedge CLK)
      state[12] <= _169_;
  always @(posedge CLK)
      state[13] <= _170_;
  always @(posedge CLK)
      state[14] <= _135_;
  always @(posedge CLK)
      state[15] <= _151_;
  always @(posedge CLK)
      state[16] <= _159_;
  always @(posedge CLK)
      state[17] <= _152_;
  always @(posedge CLK)
      state[18] <= _160_;
  always @(posedge CLK)
      state[19] <= _161_;
  always @(posedge CLK)
      state[20] <= _153_;
  always @(posedge CLK)
      state[21] <= _162_;
  always @(posedge CLK)
      state[22] <= _163_;
  always @(posedge CLK)
      state[23] <= _164_;
  always @(posedge CLK)
      state[24] <= _165_;
  always @(posedge CLK)
      state[25] <= _154_;
  always @(posedge CLK)
      state[26] <= _166_;
  assign GOOD = state[10];
endmodule
